
module fir_filter_control(

);

endmodule /* fir_filter_control */
