
module fir_filter();

endmodule /* fir_filter */

