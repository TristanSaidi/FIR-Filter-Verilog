
`timescale 1ns/1ps
`define QSIM_IN_FN_1 		"./reports/golden_block.rpt"
`define QSIM_OUT_FN_1		"./reports/outputs.rpt"
`define HALF_FAST_CLK_CYCLE	#2.00
`define HALF_SLOW_CLK_CYCLE	#20.00
`define FAST_SLOW_CLK_RATIO	10
`define QRTR_FAST_CLK_CYCLE	#1.00
`define QRTR_SLOW_CLK_CYCLE	#10.00
`define ITER 			10
`define PRECOMP			2048

module testbench();

	integer	qsim_in_1, qsim_out_1;
	integer	i;
	integer	writing;


	wire	[15:0]		Y;
	wire			valid_out;
	reg	[15:0]		X;
	reg	[19:0]		CIN;
	reg	[10:0]		CADDR;
	reg			CLOAD;
	reg			valid_in;
	reg			clk_slow, clk_fast;
	reg			resetn;
	integer 		COEF_ARRAY		[63:0];
	integer 		COMP_ARRAY		[63:0];
	integer 		COUNT_REG;
	integer	CIN_INT;
	integer	X_INT;
	integer	Y_INT;
	integer k;

	fir_filter	DUT(
		.dout		(Y),
		.valid_out	(valid_out),
		.din		(X),
		.CIN		(CIN),
		.CADDR		(CADDR),
		.CLOAD		(CLOAD),
		.valid_in	(valid_in),
		.clk_fast	(clk_fast),
		.clk_slow	(clk_slow),
		.resetn		(resetn)
	);

	always begin
		`HALF_FAST_CLK_CYCLE
		clk_fast	= ~clk_fast;
	end
	always begin
		`HALF_SLOW_CLK_CYCLE;
		clk_slow	= ~clk_slow;
	end

	integer	j;
	always	@(posedge clk_fast) begin
		j = j + 1;
	end
	always	@(negedge clk_fast) begin
		`QRTR_FAST_CLK_CYCLE;
		if (((j + 1) % `FAST_SLOW_CLK_RATIO) == 0) begin
			if (writing == 1) begin
				CIN_INT		= COMP_ARRAY[i];
				CIN		= CIN_INT;
				CADDR		= i;
				$fwrite(qsim_out_1, "%0d\n", CIN_INT);

			end
			else if (writing == 0) begin
				$fwrite(qsim_out_1, "%0d,%0d\n", X_INT, Y_INT);
				X		= i;
				X_INT		= X;
			end
		end
	end

	initial begin
		writing		= 3;
		qsim_out_1	= $fopen(`QSIM_OUT_FN_1, "w");
		clk_slow	= 0;
		clk_fast	= 0;
		resetn 		= 0;
		valid_in	= 0;
		for (k = 0; k < 64; k = k+1) begin
			@(posedge clk_fast);
			COMP_ARRAY[k] = 0;
			COEF_ARRAY[k] = $urandom%65535;		
		end
		for (k = 0; k < 8; k = k+1) begin
			for (COUNT_REG = 0; COUNT_REG < 256; COUNT_REG = COUNT_REG+1) begin
				@(posedge clk_slow);
				if(COUNT_REG == 1)begin
					COMP_ARRAY[j*8] = COMP_ARRAY[j*8] + COEF_ARRAY[j*8];
				end
				if(COUNT_REG>>1 == 1)begin
					COMP_ARRAY[j*8+1] = COMP_ARRAY[j*8+1] + COEF_ARRAY[j*8+1];
				end
				if(COUNT_REG>>2 == 1)begin
					COMP_ARRAY[j*8+2] = COMP_ARRAY[j*8+2] + COEF_ARRAY[j*8+2];
				end
				if(COUNT_REG>>3 == 1)begin
					COMP_ARRAY[j*8+3] = COMP_ARRAY[j*8+3] + COEF_ARRAY[j*8+3];
				end
				if(COUNT_REG>>4 == 1)begin
					COMP_ARRAY[j*8+4] = COMP_ARRAY[j*8+4] + COEF_ARRAY[j*8+4];
				end
				if(COUNT_REG>>5 == 1)begin
					COMP_ARRAY[j*8+5] = COMP_ARRAY[j*8+5] + COEF_ARRAY[j*8+5];
				end
				if(COUNT_REG>>6 == 1)begin
					COMP_ARRAY[j*8+6] = COMP_ARRAY[j*8+6] + COEF_ARRAY[j*8+6];
				end
				if(COUNT_REG>>7 == 1)begin
					COMP_ARRAY[j*8+7] = COMP_ARRAY[j*8+7] + COEF_ARRAY[j*8+7];
				end

			end
		end
		@(posedge clk_slow);
		clk_fast	= 1;
		@(posedge clk_slow);
		resetn 		= 1;
		CLOAD		= 1;
		writing		= 1;
		j		= 0;
		for (i = 0; i < `PRECOMP; i = i + 1) begin
			@(posedge clk_slow);
		end
		CLOAD		= 0;
		valid_in 	= 1;
		resetn		= 1;
		writing		= 0;
		j		= 0;
		for (i = 0; i < `ITER; i = i + 1) begin
			@(posedge clk_slow);
		end
		$fclose(qsim_in_1);
		$fclose(qsim_out_1);
		$finish;
	end

endmodule /* testbench */

